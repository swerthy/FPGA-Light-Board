module LightBoard(
	input CLOCK_50,
	input [3:0]KEY,
	input [9:0]SW,
	output [9:0]LEDR
	);
	
	wire clk;
	assign clk = CLOCK_50;
	wire rst;
	assign rst = KEY[0];
	wire send;
	assign send = !KEY[1];
	wire enter;
	assign enter = !KEY[3];
	wire [5642:0]bo;
	assign bo = 5643'b11000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000111000000001110000000011100000000100000000000;
	reg [5642:0]data;
	reg shifted;
	wire out;
	wire done;
 
	reg [8:0]addr;
	reg [7:0]val;
	reg [2:0]q;
	reg [4:0]qstack;
	assign LEDR[4:0] = qstack;
	
	reg [5642:0]q0;
	reg [9:0]t0;	
	
	reg [5642:0]q1;
	reg [9:0]t1;
	
	reg [5642:0]q2;
	reg [9:0]t2;
	
	reg [5642:0]q3;
	reg [9:0]t3;
	
	reg [5642:0]q4;
	reg [9:0]t4;
	
	reg [4:0]S;
	reg [4:0]NS;
	
	assign LEDR[9:5] = S;
	
	parameter 
		HOME=5'd0, 		//Home
		//Modify Address (val[1:0]==2'b11)
		ADDRX=5'd1, 	//Address selection debounce
		ADDR=5'd2, 		//Address selection
		VALX=5'd3,		//Value selection debounce
		VAL=5'd4,		//Value selection
		RECAX=5'd5,		//Record address debounce
		RECA=5'd6,		//Record address
		//Modify Cue (val[1:0]==2'b10)
		QNUMX=5'd7,		//Cue selection debounce
		QNUM=5'd8,		//Cue selection
		TIMEX=5'd9,		//Fade time selection debounce
		TIME=5'd10,		//Fade time selection
		RECQX=5'd11,	//Record cue debounce
		RECQ=5'd12,		//Record cue
		//Go to Cue (val[1:0]==2'b01)
		QGOX=5'd13,		//Destination selection debounce
		QGO=5'd14,		//Destination selection
		SETX=5'd15,		//Set cue debounce
		SET=5'd16,		//Set cue
		//Go to next cue (val[1:0]==2'b00)
		SHIFT=5'd17,	//Fade
		//Other
		ERROR=5'hff;
		
		
	always@(posedge clk or negedge rst)
		if(rst==1'b0)
			S <= HOME;
		else
			S <= NS;

	always@(*)
		case(S)
			
			HOME:
			begin
				if(enter==0)
					NS <= HOME;
				else
				begin
					case(SW[1:0])
						
						2'b11: NS <= ADDRX;
						2'b10: NS <= QNUMX;
						2'b01: NS <= QGOX;
						2'b00: NS <= SHIFT;
						
					endcase
				end
			end
			
			ADDRX: 
			if(enter==1)
				NS <= ADDRX;
			else
				NS <= ADDR;
			
			ADDR:
			if(enter==0)
				NS <= ADDR;
			else
				NS <= VALX;
			
			VALX:
			if(enter==1)
				NS <= VALX;
			else
				NS <= VAL;
			
			VAL:
			if(enter==0)
				NS <= VAL;
			else
				NS <= RECAX;
			
			RECAX:
			if(enter==1)
				NS <= RECAX;
			else
				NS <= RECA;
				
			RECA: NS <= HOME;
			
			QNUMX:
			if(enter==1)
				NS <= QNUMX;
			else
				NS <= QNUM;
				
			QNUM:
			if(enter==0)
				NS <= QNUM;
			else
				NS <= TIMEX;
			
			TIMEX:
			if(enter==1)
				NS <= TIMEX;
			else
				NS <= TIME;
			
			TIME:
			if(enter==0)
				NS <= TIME;
			else
				NS <= RECQX;
			
			RECQX:
			if(enter==1)
				NS <= RECQX;
			else
				NS <= RECQ;
			
			RECQ: NS <= HOME;
			
			QGOX:
			if(enter==1)
				NS <= QGOX;
			else
				NS <= QGO;
			
			QGO:
			if(enter==0)
				NS <= QGO;
			else
				NS <= SETX;
			
			SETX:
			if(enter==1)
				NS <= SETX;
			else
				NS <= SET;
			
			SET: NS <= HOME;
			
			SHIFT:
			if(shifted==1)
				NS <= HOME;
			else
				NS <= SHIFT;

		endcase

	always@(posedge clk or negedge rst)
		if(rst==1'b0)
		begin
			data <= bo;
			q0 <= bo;
			q1 <= bo;
			q2 <= bo;
			q3 <= bo;
			q4 <= bo;
			t0 <= 10'd0;
			t1 <= 10'd0;
			t2 <= 10'd0;
			t3 <= 10'd0;
			t4 <= 10'd0;	
			qstack <= 5'b00000;
		end
		else
		begin
		case(S)
			
//			HOME: 
		
			ADDRX: addr <= SW[8:0];
			
			ADDR: addr <= SW[8:0];
			
			VALX: val <= SW[7:0];

			VAL: val <= SW[7:0]; 
			
			RECAX: 
			
			RECA: 
			case(addr)
				9'd1: val <= [12:19];
				9'd2: val <= [23:30];
				9'd3: val <= [34:41];
				9'd4: val <= [45:52];
				9'd5: val <= [56:63];
				9'd6: val <= [67:74];
				9'd7: val <= [78:85];
				9'd8: val <= [89:96];
				9'd9: val <= [100:107];
				9'd10: val <= [111:118];
				9'd11: val <= [122:129];
				9'd12: val <= [133:140];
				9'd13: val <= [144:151];
				9'd14: val <= [155:162];
				9'd15: val <= [166:173];
				9'd16: val <= [177:184];
				9'd17: val <= [188:195];
				9'd18: val <= [199:206];
				9'd19: val <= [210:217];
				9'd20: val <= [221:228];
				9'd21: val <= [232:239];
				9'd22: val <= [243:250];
				9'd23: val <= [254:261];
				9'd24: val <= [265:272];
				9'd25: val <= [276:283];
				9'd26: val <= [287:294];
				9'd27: val <= [298:305];
				9'd28: val <= [309:316];
				9'd29: val <= [320:327];
				9'd30: val <= [331:338];
				9'd31: val <= [342:349];
				9'd32: val <= [353:360];
				9'd33: val <= [364:371];
				9'd34: val <= [375:382];
				9'd35: val <= [386:393];
				9'd36: val <= [397:404];
				9'd37: val <= [408:415];
				9'd38: val <= [419:426];
				9'd39: val <= [430:437];
				9'd40: val <= [441:448];
				9'd41: val <= [452:459];
				9'd42: val <= [463:470];
				9'd43: val <= [474:481];
				9'd44: val <= [485:492];
				9'd45: val <= [496:503];
				9'd46: val <= [507:514];
				9'd47: val <= [518:525];
				9'd48: val <= [529:536];
				9'd49: val <= [540:547];
				9'd50: val <= [551:558];
				9'd51: val <= [562:569];
				9'd52: val <= [573:580];
				9'd53: val <= [584:591];
				9'd54: val <= [595:602];
				9'd55: val <= [606:613];
				9'd56: val <= [617:624];
				9'd57: val <= [628:635];
				9'd58: val <= [639:646];
				9'd59: val <= [650:657];
				9'd60: val <= [661:668];
				9'd61: val <= [672:679];
				9'd62: val <= [683:690];
				9'd63: val <= [694:701];
				9'd64: val <= [705:712];
				9'd65: val <= [716:723];
				9'd66: val <= [727:734];
				9'd67: val <= [738:745];
				9'd68: val <= [749:756];
				9'd69: val <= [760:767];
				9'd70: val <= [771:778];
				9'd71: val <= [782:789];
				9'd72: val <= [793:800];
				9'd73: val <= [804:811];
				9'd74: val <= [815:822];
				9'd75: val <= [826:833];
				9'd76: val <= [837:844];
				9'd77: val <= [848:855];
				9'd78: val <= [859:866];
				9'd79: val <= [870:877];
				9'd80: val <= [881:888];
				9'd81: val <= [892:899];
				9'd82: val <= [903:910];
				9'd83: val <= [914:921];
				9'd84: val <= [925:932];
				9'd85: val <= [936:943];
				9'd86: val <= [947:954];
				9'd87: val <= [958:965];
				9'd88: val <= [969:976];
				9'd89: val <= [980:987];
				9'd90: val <= [991:998];
				9'd91: val <= [1002:1009];
				9'd92: val <= [1013:1020];
				9'd93: val <= [1024:1031];
				9'd94: val <= [1035:1042];
				9'd95: val <= [1046:1053];
				9'd96: val <= [1057:1064];
				9'd97: val <= [1068:1075];
				9'd98: val <= [1079:1086];
				9'd99: val <= [1090:1097];
				9'd100: val <= [1101:1108];
				9'd101: val <= [1112:1119];
				9'd102: val <= [1123:1130];
				9'd103: val <= [1134:1141];
				9'd104: val <= [1145:1152];
				9'd105: val <= [1156:1163];
				9'd106: val <= [1167:1174];
				9'd107: val <= [1178:1185];
				9'd108: val <= [1189:1196];
				9'd109: val <= [1200:1207];
				9'd110: val <= [1211:1218];
				9'd111: val <= [1222:1229];
				9'd112: val <= [1233:1240];
				9'd113: val <= [1244:1251];
				9'd114: val <= [1255:1262];
				9'd115: val <= [1266:1273];
				9'd116: val <= [1277:1284];
				9'd117: val <= [1288:1295];
				9'd118: val <= [1299:1306];
				9'd119: val <= [1310:1317];
				9'd120: val <= [1321:1328];
				9'd121: val <= [1332:1339];
				9'd122: val <= [1343:1350];
				9'd123: val <= [1354:1361];
				9'd124: val <= [1365:1372];
				9'd125: val <= [1376:1383];
				9'd126: val <= [1387:1394];
				9'd127: val <= [1398:1405];
				9'd128: val <= [1409:1416];
				9'd129: val <= [1420:1427];
				9'd130: val <= [1431:1438];
				9'd131: val <= [1442:1449];
				9'd132: val <= [1453:1460];
				9'd133: val <= [1464:1471];
				9'd134: val <= [1475:1482];
				9'd135: val <= [1486:1493];
				9'd136: val <= [1497:1504];
				9'd137: val <= [1508:1515];
				9'd138: val <= [1519:1526];
				9'd139: val <= [1530:1537];
				9'd140: val <= [1541:1548];
				9'd141: val <= [1552:1559];
				9'd142: val <= [1563:1570];
				9'd143: val <= [1574:1581];
				9'd144: val <= [1585:1592];
				9'd145: val <= [1596:1603];
				9'd146: val <= [1607:1614];
				9'd147: val <= [1618:1625];
				9'd148: val <= [1629:1636];
				9'd149: val <= [1640:1647];
				9'd150: val <= [1651:1658];
				9'd151: val <= [1662:1669];
				9'd152: val <= [1673:1680];
				9'd153: val <= [1684:1691];
				9'd154: val <= [1695:1702];
				9'd155: val <= [1706:1713];
				9'd156: val <= [1717:1724];
				9'd157: val <= [1728:1735];
				9'd158: val <= [1739:1746];
				9'd159: val <= [1750:1757];
				9'd160: val <= [1761:1768];
				9'd161: val <= [1772:1779];
				9'd162: val <= [1783:1790];
				9'd163: val <= [1794:1801];
				9'd164: val <= [1805:1812];
				9'd165: val <= [1816:1823];
				9'd166: val <= [1827:1834];
				9'd167: val <= [1838:1845];
				9'd168: val <= [1849:1856];
				9'd169: val <= [1860:1867];
				9'd170: val <= [1871:1878];
				9'd171: val <= [1882:1889];
				9'd172: val <= [1893:1900];
				9'd173: val <= [1904:1911];
				9'd174: val <= [1915:1922];
				9'd175: val <= [1926:1933];
				9'd176: val <= [1937:1944];
				9'd177: val <= [1948:1955];
				9'd178: val <= [1959:1966];
				9'd179: val <= [1970:1977];
				9'd180: val <= [1981:1988];
				9'd181: val <= [1992:1999];
				9'd182: val <= [2003:2010];
				9'd183: val <= [2014:2021];
				9'd184: val <= [2025:2032];
				9'd185: val <= [2036:2043];
				9'd186: val <= [2047:2054];
				9'd187: val <= [2058:2065];
				9'd188: val <= [2069:2076];
				9'd189: val <= [2080:2087];
				9'd190: val <= [2091:2098];
				9'd191: val <= [2102:2109];
				9'd192: val <= [2113:2120];
				9'd193: val <= [2124:2131];
				9'd194: val <= [2135:2142];
				9'd195: val <= [2146:2153];
				9'd196: val <= [2157:2164];
				9'd197: val <= [2168:2175];
				9'd198: val <= [2179:2186];
				9'd199: val <= [2190:2197];
				9'd200: val <= [2201:2208];
				9'd201: val <= [2212:2219];
				9'd202: val <= [2223:2230];
				9'd203: val <= [2234:2241];
				9'd204: val <= [2245:2252];
				9'd205: val <= [2256:2263];
				9'd206: val <= [2267:2274];
				9'd207: val <= [2278:2285];
				9'd208: val <= [2289:2296];
				9'd209: val <= [2300:2307];
				9'd210: val <= [2311:2318];
				9'd211: val <= [2322:2329];
				9'd212: val <= [2333:2340];
				9'd213: val <= [2344:2351];
				9'd214: val <= [2355:2362];
				9'd215: val <= [2366:2373];
				9'd216: val <= [2377:2384];
				9'd217: val <= [2388:2395];
				9'd218: val <= [2399:2406];
				9'd219: val <= [2410:2417];
				9'd220: val <= [2421:2428];
				9'd221: val <= [2432:2439];
				9'd222: val <= [2443:2450];
				9'd223: val <= [2454:2461];
				9'd224: val <= [2465:2472];
				9'd225: val <= [2476:2483];
				9'd226: val <= [2487:2494];
				9'd227: val <= [2498:2505];
				9'd228: val <= [2509:2516];
				9'd229: val <= [2520:2527];
				9'd230: val <= [2531:2538];
				9'd231: val <= [2542:2549];
				9'd232: val <= [2553:2560];
				9'd233: val <= [2564:2571];
				9'd234: val <= [2575:2582];
				9'd235: val <= [2586:2593];
				9'd236: val <= [2597:2604];
				9'd237: val <= [2608:2615];
				9'd238: val <= [2619:2626];
				9'd239: val <= [2630:2637];
				9'd240: val <= [2641:2648];
				9'd241: val <= [2652:2659];
				9'd242: val <= [2663:2670];
				9'd243: val <= [2674:2681];
				9'd244: val <= [2685:2692];
				9'd245: val <= [2696:2703];
				9'd246: val <= [2707:2714];
				9'd247: val <= [2718:2725];
				9'd248: val <= [2729:2736];
				9'd249: val <= [2740:2747];
				9'd250: val <= [2751:2758];
				9'd251: val <= [2762:2769];
				9'd252: val <= [2773:2780];
				9'd253: val <= [2784:2791];
				9'd254: val <= [2795:2802];
				9'd255: val <= [2806:2813];
				9'd256: val <= [2817:2824];
				9'd257: val <= [2828:2835];
				9'd258: val <= [2839:2846];
				9'd259: val <= [2850:2857];
				9'd260: val <= [2861:2868];
				9'd261: val <= [2872:2879];
				9'd262: val <= [2883:2890];
				9'd263: val <= [2894:2901];
				9'd264: val <= [2905:2912];
				9'd265: val <= [2916:2923];
				9'd266: val <= [2927:2934];
				9'd267: val <= [2938:2945];
				9'd268: val <= [2949:2956];
				9'd269: val <= [2960:2967];
				9'd270: val <= [2971:2978];
				9'd271: val <= [2982:2989];
				9'd272: val <= [2993:3000];
				9'd273: val <= [3004:3011];
				9'd274: val <= [3015:3022];
				9'd275: val <= [3026:3033];
				9'd276: val <= [3037:3044];
				9'd277: val <= [3048:3055];
				9'd278: val <= [3059:3066];
				9'd279: val <= [3070:3077];
				9'd280: val <= [3081:3088];
				9'd281: val <= [3092:3099];
				9'd282: val <= [3103:3110];
				9'd283: val <= [3114:3121];
				9'd284: val <= [3125:3132];
				9'd285: val <= [3136:3143];
				9'd286: val <= [3147:3154];
				9'd287: val <= [3158:3165];
				9'd288: val <= [3169:3176];
				9'd289: val <= [3180:3187];
				9'd290: val <= [3191:3198];
				9'd291: val <= [3202:3209];
				9'd292: val <= [3213:3220];
				9'd293: val <= [3224:3231];
				9'd294: val <= [3235:3242];
				9'd295: val <= [3246:3253];
				9'd296: val <= [3257:3264];
				9'd297: val <= [3268:3275];
				9'd298: val <= [3279:3286];
				9'd299: val <= [3290:3297];
				9'd300: val <= [3301:3308];
				9'd301: val <= [3312:3319];
				9'd302: val <= [3323:3330];
				9'd303: val <= [3334:3341];
				9'd304: val <= [3345:3352];
				9'd305: val <= [3356:3363];
				9'd306: val <= [3367:3374];
				9'd307: val <= [3378:3385];
				9'd308: val <= [3389:3396];
				9'd309: val <= [3400:3407];
				9'd310: val <= [3411:3418];
				9'd311: val <= [3422:3429];
				9'd312: val <= [3433:3440];
				9'd313: val <= [3444:3451];
				9'd314: val <= [3455:3462];
				9'd315: val <= [3466:3473];
				9'd316: val <= [3477:3484];
				9'd317: val <= [3488:3495];
				9'd318: val <= [3499:3506];
				9'd319: val <= [3510:3517];
				9'd320: val <= [3521:3528];
				9'd321: val <= [3532:3539];
				9'd322: val <= [3543:3550];
				9'd323: val <= [3554:3561];
				9'd324: val <= [3565:3572];
				9'd325: val <= [3576:3583];
				9'd326: val <= [3587:3594];
				9'd327: val <= [3598:3605];
				9'd328: val <= [3609:3616];
				9'd329: val <= [3620:3627];
				9'd330: val <= [3631:3638];
				9'd331: val <= [3642:3649];
				9'd332: val <= [3653:3660];
				9'd333: val <= [3664:3671];
				9'd334: val <= [3675:3682];
				9'd335: val <= [3686:3693];
				9'd336: val <= [3697:3704];
				9'd337: val <= [3708:3715];
				9'd338: val <= [3719:3726];
				9'd339: val <= [3730:3737];
				9'd340: val <= [3741:3748];
				9'd341: val <= [3752:3759];
				9'd342: val <= [3763:3770];
				9'd343: val <= [3774:3781];
				9'd344: val <= [3785:3792];
				9'd345: val <= [3796:3803];
				9'd346: val <= [3807:3814];
				9'd347: val <= [3818:3825];
				9'd348: val <= [3829:3836];
				9'd349: val <= [3840:3847];
				9'd350: val <= [3851:3858];
				9'd351: val <= [3862:3869];
				9'd352: val <= [3873:3880];
				9'd353: val <= [3884:3891];
				9'd354: val <= [3895:3902];
				9'd355: val <= [3906:3913];
				9'd356: val <= [3917:3924];
				9'd357: val <= [3928:3935];
				9'd358: val <= [3939:3946];
				9'd359: val <= [3950:3957];
				9'd360: val <= [3961:3968];
				9'd361: val <= [3972:3979];
				9'd362: val <= [3983:3990];
				9'd363: val <= [3994:4001];
				9'd364: val <= [4005:4012];
				9'd365: val <= [4016:4023];
				9'd366: val <= [4027:4034];
				9'd367: val <= [4038:4045];
				9'd368: val <= [4049:4056];
				9'd369: val <= [4060:4067];
				9'd370: val <= [4071:4078];
				9'd371: val <= [4082:4089];
				9'd372: val <= [4093:4100];
				9'd373: val <= [4104:4111];
				9'd374: val <= [4115:4122];
				9'd375: val <= [4126:4133];
				9'd376: val <= [4137:4144];
				9'd377: val <= [4148:4155];
				9'd378: val <= [4159:4166];
				9'd379: val <= [4170:4177];
				9'd380: val <= [4181:4188];
				9'd381: val <= [4192:4199];
				9'd382: val <= [4203:4210];
				9'd383: val <= [4214:4221];
				9'd384: val <= [4225:4232];
				9'd385: val <= [4236:4243];
				9'd386: val <= [4247:4254];
				9'd387: val <= [4258:4265];
				9'd388: val <= [4269:4276];
				9'd389: val <= [4280:4287];
				9'd390: val <= [4291:4298];
				9'd391: val <= [4302:4309];
				9'd392: val <= [4313:4320];
				9'd393: val <= [4324:4331];
				9'd394: val <= [4335:4342];
				9'd395: val <= [4346:4353];
				9'd396: val <= [4357:4364];
				9'd397: val <= [4368:4375];
				9'd398: val <= [4379:4386];
				9'd399: val <= [4390:4397];
				9'd400: val <= [4401:4408];
				9'd401: val <= [4412:4419];
				9'd402: val <= [4423:4430];
				9'd403: val <= [4434:4441];
				9'd404: val <= [4445:4452];
				9'd405: val <= [4456:4463];
				9'd406: val <= [4467:4474];
				9'd407: val <= [4478:4485];
				9'd408: val <= [4489:4496];
				9'd409: val <= [4500:4507];
				9'd410: val <= [4511:4518];
				9'd411: val <= [4522:4529];
				9'd412: val <= [4533:4540];
				9'd413: val <= [4544:4551];
				9'd414: val <= [4555:4562];
				9'd415: val <= [4566:4573];
				9'd416: val <= [4577:4584];
				9'd417: val <= [4588:4595];
				9'd418: val <= [4599:4606];
				9'd419: val <= [4610:4617];
				9'd420: val <= [4621:4628];
				9'd421: val <= [4632:4639];
				9'd422: val <= [4643:4650];
				9'd423: val <= [4654:4661];
				9'd424: val <= [4665:4672];
				9'd425: val <= [4676:4683];
				9'd426: val <= [4687:4694];
				9'd427: val <= [4698:4705];
				9'd428: val <= [4709:4716];
				9'd429: val <= [4720:4727];
				9'd430: val <= [4731:4738];
				9'd431: val <= [4742:4749];
				9'd432: val <= [4753:4760];
				9'd433: val <= [4764:4771];
				9'd434: val <= [4775:4782];
				9'd435: val <= [4786:4793];
				9'd436: val <= [4797:4804];
				9'd437: val <= [4808:4815];
				9'd438: val <= [4819:4826];
				9'd439: val <= [4830:4837];
				9'd440: val <= [4841:4848];
				9'd441: val <= [4852:4859];
				9'd442: val <= [4863:4870];
				9'd443: val <= [4874:4881];
				9'd444: val <= [4885:4892];
				9'd445: val <= [4896:4903];
				9'd446: val <= [4907:4914];
				9'd447: val <= [4918:4925];
				9'd448: val <= [4929:4936];
				9'd449: val <= [4940:4947];
				9'd450: val <= [4951:4958];
				9'd451: val <= [4962:4969];
				9'd452: val <= [4973:4980];
				9'd453: val <= [4984:4991];
				9'd454: val <= [4995:5002];
				9'd455: val <= [5006:5013];
				9'd456: val <= [5017:5024];
				9'd457: val <= [5028:5035];
				9'd458: val <= [5039:5046];
				9'd459: val <= [5050:5057];
				9'd460: val <= [5061:5068];
				9'd461: val <= [5072:5079];
				9'd462: val <= [5083:5090];
				9'd463: val <= [5094:5101];
				9'd464: val <= [5105:5112];
				9'd465: val <= [5116:5123];
				9'd466: val <= [5127:5134];
				9'd467: val <= [5138:5145];
				9'd468: val <= [5149:5156];
				9'd469: val <= [5160:5167];
				9'd470: val <= [5171:5178];
				9'd471: val <= [5182:5189];
				9'd472: val <= [5193:5200];
				9'd473: val <= [5204:5211];
				9'd474: val <= [5215:5222];
				9'd475: val <= [5226:5233];
				9'd476: val <= [5237:5244];
				9'd477: val <= [5248:5255];
				9'd478: val <= [5259:5266];
				9'd479: val <= [5270:5277];
				9'd480: val <= [5281:5288];
				9'd481: val <= [5292:5299];
				9'd482: val <= [5303:5310];
				9'd483: val <= [5314:5321];
				9'd484: val <= [5325:5332];
				9'd485: val <= [5336:5343];
				9'd486: val <= [5347:5354];
				9'd487: val <= [5358:5365];
				9'd488: val <= [5369:5376];
				9'd489: val <= [5380:5387];
				9'd490: val <= [5391:5398];
				9'd491: val <= [5402:5409];
				9'd492: val <= [5413:5420];
				9'd493: val <= [5424:5431];
				9'd494: val <= [5435:5442];
				9'd495: val <= [5446:5453];
				9'd496: val <= [5457:5464];
				9'd497: val <= [5468:5475];
				9'd498: val <= [5479:5486];
				9'd499: val <= [5490:5497];
				9'd500: val <= [5501:5508];
				9'd501: val <= [5512:5519];
				9'd502: val <= [5523:5530];
				9'd503: val <= [5534:5541];
				9'd504: val <= [5545:5552];
				9'd505: val <= [5556:5563];
				9'd506: val <= [5567:5574];
				9'd507: val <= [5578:5585];
				9'd508: val <= [5589:5596];
				9'd509: val <= [5600:5607];
				9'd510: val <= [5611:5618];
				9'd511: val <= [5622:5629];
			endcase
			
			QNUMX: q <= SW[2:0];
			
			QNUM: q <= SW[2:0];
			
			TIMEX: 
			case(q)
				3'd0: t0 <= SW[9:0];
				3'd1: t1 <= SW[9:0];
				3'd2: t2 <= SW[9:0];
				3'd3: t3 <= SW[9:0];
				3'd4: t4 <= SW[9:0];
//				default: S <= ERROR;
			endcase
			
			TIME:
			case(q)
				3'd0: t0 <= SW[9:0];
				3'd1: t1 <= SW[9:0];
				3'd2: t2 <= SW[9:0];
				3'd3: t3 <= SW[9:0];
				3'd4: t4 <= SW[9:0];
//				default: S <= ERROR;
			endcase
			
			RECQX:
			case(q)
			
				3'd0: 
				begin
					q0 <= data;
					qstack[0] <= 1;
				end
				
				3'd1: 
				begin
					q1 <= data;
					qstack[1] <= 1;
				end
				
				3'd2: 
				begin
					q2 <= data;
					qstack[2] <= 1;
				end
				
				3'd3: 
				begin
					q3 <= data;
					qstack[3] <= 1;
				end
				
				3'd4: 
				begin
					q4 <= data;
					qstack[4] <= 1;
				end
				
//				default: S <= ERROR;
				
			endcase
			
			RECQ:
			case(q)
			
				3'd0: 
				begin
					q0 <= data;
					qstack[0] <= 1;
				end
				
				3'd1: 
				begin
					q1 <= data;
					qstack[1] <= 1;
				end
				
				3'd2: 
				begin
					q2 <= data;
					qstack[2] <= 1;
				end
				
				3'd3: 
				begin
					q3 <= data;
					qstack[3] <= 1;
				end
				
				3'd4: 
				begin
					q4 <= data;
					qstack[4] <= 1;
				end
				
//				default: S <= ERROR;
				
			endcase
			
			QGOX: q <= SW[2:0];
			
			QGO: q <= SW[2:0];
			
			SETX: 
			case(q)
				3'd0: data <= q0;
				3'd1: data <= q1;
				3'd2: data <= q2;
				3'd3: data <= q3;
				3'd4: data <= q4;
//				default: S <= ERROR;
			endcase
			
			SET: 
			case(q)
				3'd0: data <= q0;
				3'd1: data <= q1;
				3'd2: data <= q2;
				3'd3: data <= q3;
				3'd4: data <= q4;
//				default: S <= ERROR;
			endcase
			
//			SHIFT:
			
		endcase
		end
	
	packet sendpacket(clk,rst,send,data,out,done);
	//packet sendpacket(clk,rst,send,data,output,done);
	
endmodule
